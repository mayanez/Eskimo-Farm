/*
 * Avalon memory-mapped peripheral for the VGA LED Emulator
 *
 * Stephen A. Edwards
 * Columbia University
 */

module VGA_LED(input logic        clk,
	       input logic 	  reset,
	       input logic [511:0] gl_input, /* 20 * 24-bit entries rounded up to closest power of 2 */
	       input logic 	  write,
	       output logic [7:0] VGA_R, VGA_G, VGA_B,
	       output logic 	  VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK_n,
	       output logic 	  VGA_SYNC_n);

   logic [23:0] gl_array [20:0];
   logic [23:0] sprite1,sprite2,sprite3,sprite4,sprite5,sprite6,sprite7,sprite8,sprite9,sprite10,sprite11,sprite12,sprite13,sprite14,sprite15,sprite16,sprite17,sprite18,sprite19,sprite20;
   logic [4:0] id1,id2,id3,id4,id5,id6,id7,id8,id9,id10,id11,id12,id13,id14,id15,id16,id17,id18,id19,id20;

   logic [9:0] VGA_HCOUNT;
   logic [9:0] VGA_VCOUNT;
   logic VGA_CLOCK;

   assign gl_array[0] = gl_input[23:0];
   assign gl_array[1] = gl_input[45:24];
   assign gl_array[2] = gl_input[68:46];
   assign gl_array[3] = gl_input[91:69];
   assign gl_array[4] = gl_input[114:92];
   assign gl_array[5] = gl_input[137:115];
   assign gl_array[6] = gl_input[160:138];
   assign gl_array[7] = gl_input[183:161];
   assign gl_array[8] = gl_input[206:184];
   assign gl_array[9] = gl_input[229:207];
   assign gl_array[10] = gl_input[252:230];
   assign gl_array[11] = gl_input[275:253];
   assign gl_array[12] = gl_input[298:276];
   assign gl_array[13] = gl_input[321:299];
   assign gl_array[14] = gl_input[344:322];
   assign gl_array[15] = gl_input[367:345];
   assign gl_array[16] = gl_input[390:368];
   assign gl_array[17] = gl_input[413:391];
   assign gl_array[18] = gl_input[436:414];
   assign gl_array[19] = gl_input[459:437];
   assign gl_array[20] = gl_input[482:460];
   assign gl_array[21] = gl_input[506:483];


   assign sprite1 = gl_array[0];
   assign sprite2 = gl_array[1];
   assign sprite3 = gl_array[2];
   assign sprite4 = gl_array[3];
   assign sprite5 = gl_array[4];
   assign sprite6 = gl_array[5];
   assign sprite7 = gl_array[6];
   assign sprite8 = gl_array[7];
   assign sprite9 = gl_array[8];
   assign sprite10 = gl_array[9];
   assign sprite11 = gl_array[10];
   assign sprite12 = gl_array[11];
   assign sprite13 = gl_array[12];
   assign sprite14 = gl_array[13];
   assign sprite15 = gl_array[14];
   assign sprite16 = gl_array[15];
   assign sprite17 = gl_array[16];
   assign sprite18 = gl_array[17];
   assign sprite19 = gl_array[18];
   assign sprite20 = gl_array[19];
   assign sprite21 = gl_array[20];

   assign id1 = sprite1[23:19];
   assign id2 = sprite2[23:19];
   assign id3 = sprite3[23:19];
   assign id4 = sprite4[23:19];
   assign id5 = sprite5[23:19];
   assign id6 = sprite6[23:19];
   assign id7 = sprite7[23:19];
   assign id8 = sprite8[23:19];
   assign id9 = sprite9[23:19];
   assign id10 = sprite10[23:19];
   assign id11 = sprite11[23:19];
   assign id12 = sprite12[23:19];
   assign id13 = sprite13[23:19];
   assign id14 = sprite14[23:19];
   assign id15 = sprite15[23:19];
   assign id16 = sprite16[23:19];
   assign id17 = sprite17[23:19];
   assign id18 = sprite18[23:19];
   assign id19 = sprite19[23:19];
   assign id20 = sprite20[23:19];
   assign id21 = sprite21[23:19];

   logic [11:0] addr_ship,addr_pig,addr_bee,addr_sheep,addr_cow,addr_hen,addr_mcdonald,addr_h_eskimo,addr_s_eskimo,addr_score,addr_one,addr_two,addr_three,addr_four,addr_five,addr_six,addr_seven,addr_eight,addr_nine,addr_zero,addr_bullet;

   logic [23:0] M_sprite1,M_sprite2,M_sprite3,M_sprite4,M_sprite5,M_sprite6,M_sprite7,M_sprite8,M_sprite9,M_sprite10,M_sprite11,M_sprite12,M_sprite13,M_sprite14,M_sprite15,M_sprite16,M_sprite17,M_sprite18,M_sprite19,M_sprite20,M_sprite21;
   
   
   assign M_sprite1 = (id1 == 5'd1) ? M_ship : 0;
   assign M_sprite1 = (id1 == 5'd2) ? M_pig : 0;
   assign M_sprite1 = (id1 == 5'd3) ? M_bee : 0;
   assign M_sprite1 = (id1 == 5'd4) ? M_sheep : 0;
   assign M_sprite1 = (id1 == 5'd5) ? M_cow : 0;
   assign M_sprite1 = (id1 == 5'd6) ? M_hen : 0;
   assign M_sprite1 = (id1 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite1 = (id1 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite1 = (id1 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite1 = (id1 == 5'd10) ? M_score : 0;
   assign M_sprite1 = (id1 == 5'd11) ? M_one : 0;
   assign M_sprite1 = (id1 == 5'd12) ? M_two : 0;
   assign M_sprite1 = (id1 == 5'd13) ? M_three : 0;
   assign M_sprite1 = (id1 == 5'd14) ? M_four : 0;
   assign M_sprite1 = (id1 == 5'd15) ? M_five : 0;
   assign M_sprite1 = (id1 == 5'd16) ? M_six : 0;
   assign M_sprite1 = (id1 == 5'd17) ? M_seven : 0;
   assign M_sprite1 = (id1 == 5'd18) ? M_eight : 0;
   assign M_sprite1 = (id1 == 5'd19) ? M_nine : 0;
   assign M_sprite1 = (id1 == 5'd20) ? M_zero : 0;
   assign M_sprite1 = (id1 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite2 = (id2 == 5'd1) ? M_ship : 0;
   assign M_sprite2 = (id2 == 5'd2) ? M_pig : 0;
   assign M_sprite2 = (id2 == 5'd3) ? M_bee : 0;
   assign M_sprite2 = (id2 == 5'd4) ? M_sheep : 0;
   assign M_sprite2 = (id2 == 5'd5) ? M_cow : 0;
   assign M_sprite2 = (id2 == 5'd6) ? M_hen : 0;
   assign M_sprite2 = (id2 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite2 = (id2 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite2 = (id2 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite2 = (id2 == 5'd10) ? M_score : 0;
   assign M_sprite2 = (id2 == 5'd11) ? M_one : 0;
   assign M_sprite2 = (id2 == 5'd12) ? M_two : 0;
   assign M_sprite2 = (id2 == 5'd13) ? M_three : 0;
   assign M_sprite2 = (id2 == 5'd14) ? M_four : 0;
   assign M_sprite2 = (id2 == 5'd15) ? M_five : 0;
   assign M_sprite2 = (id2 == 5'd16) ? M_six : 0;
   assign M_sprite2 = (id2 == 5'd17) ? M_seven : 0;
   assign M_sprite2 = (id2 == 5'd18) ? M_eight : 0;
   assign M_sprite2 = (id2 == 5'd19) ? M_nine : 0;
   assign M_sprite2 = (id2 == 5'd20) ? M_zero : 0;
   assign M_sprite2 = (id2 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite3 = (id3 == 5'd1) ? M_ship : 0;
   assign M_sprite3 = (id3 == 5'd2) ? M_pig : 0;
   assign M_sprite3 = (id3 == 5'd3) ? M_bee : 0;
   assign M_sprite3 = (id3 == 5'd4) ? M_sheep : 0;
   assign M_sprite3 = (id3 == 5'd5) ? M_cow : 0;
   assign M_sprite3 = (id3 == 5'd6) ? M_hen : 0;
   assign M_sprite3 = (id3 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite3 = (id3 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite3 = (id3 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite3 = (id3 == 5'd10) ? M_score : 0;
   assign M_sprite3 = (id3 == 5'd11) ? M_one : 0;
   assign M_sprite3 = (id3 == 5'd12) ? M_two : 0;
   assign M_sprite3 = (id3 == 5'd13) ? M_three : 0;
   assign M_sprite3 = (id3 == 5'd14) ? M_four : 0;
   assign M_sprite3 = (id3 == 5'd15) ? M_five : 0;
   assign M_sprite3 = (id3 == 5'd16) ? M_six : 0;
   assign M_sprite3 = (id3 == 5'd17) ? M_seven : 0;
   assign M_sprite3 = (id3 == 5'd18) ? M_eight : 0;
   assign M_sprite3 = (id3 == 5'd19) ? M_nine : 0;
   assign M_sprite3 = (id3 == 5'd20) ? M_zero : 0;
   assign M_sprite3 = (id3 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite4 = (id4 == 5'd1) ? M_ship : 0;
   assign M_sprite4 = (id4 == 5'd2) ? M_pig : 0;
   assign M_sprite4 = (id4 == 5'd3) ? M_bee : 0;
   assign M_sprite4 = (id4 == 5'd4) ? M_sheep : 0;
   assign M_sprite4 = (id4 == 5'd5) ? M_cow : 0;
   assign M_sprite4 = (id4 == 5'd6) ? M_hen : 0;
   assign M_sprite4 = (id4 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite4 = (id4 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite4 = (id4 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite4 = (id4 == 5'd10) ? M_score : 0;
   assign M_sprite4 = (id4 == 5'd11) ? M_one : 0;
   assign M_sprite4 = (id4 == 5'd12) ? M_two : 0;
   assign M_sprite4 = (id4 == 5'd13) ? M_three : 0;
   assign M_sprite4 = (id4 == 5'd14) ? M_four : 0;
   assign M_sprite4 = (id4 == 5'd15) ? M_five : 0;
   assign M_sprite4 = (id4 == 5'd16) ? M_six : 0;
   assign M_sprite4 = (id4 == 5'd17) ? M_seven : 0;
   assign M_sprite4 = (id4 == 5'd18) ? M_eight : 0;
   assign M_sprite4 = (id4 == 5'd19) ? M_nine : 0;
   assign M_sprite4 = (id4 == 5'd20) ? M_zero : 0;
   assign M_sprite4 = (id4 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite5 = (id5 == 5'd1) ? M_ship : 0;
   assign M_sprite5 = (id5 == 5'd2) ? M_pig : 0;
   assign M_sprite5 = (id5 == 5'd3) ? M_bee : 0;
   assign M_sprite5 = (id5 == 5'd4) ? M_sheep : 0;
   assign M_sprite5 = (id5 == 5'd5) ? M_cow : 0;
   assign M_sprite5 = (id5 == 5'd6) ? M_hen : 0;
   assign M_sprite5 = (id5 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite5 = (id5 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite5 = (id5 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite5 = (id5 == 5'd10) ? M_score : 0;
   assign M_sprite5 = (id5 == 5'd11) ? M_one : 0;
   assign M_sprite5 = (id5 == 5'd12) ? M_two : 0;
   assign M_sprite5 = (id5 == 5'd13) ? M_three : 0;
   assign M_sprite5 = (id5 == 5'd14) ? M_four : 0;
   assign M_sprite5 = (id5 == 5'd15) ? M_five : 0;
   assign M_sprite5 = (id5 == 5'd16) ? M_six : 0;
   assign M_sprite5 = (id5 == 5'd17) ? M_seven : 0;
   assign M_sprite5 = (id5 == 5'd18) ? M_eight : 0;
   assign M_sprite5 = (id5 == 5'd19) ? M_nine : 0;
   assign M_sprite5 = (id5 == 5'd20) ? M_zero : 0;
   assign M_sprite5 = (id5 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite6 = (id6 == 5'd1) ? M_ship : 0;
   assign M_sprite6 = (id6 == 5'd2) ? M_pig : 0;
   assign M_sprite6 = (id6 == 5'd3) ? M_bee : 0;
   assign M_sprite6 = (id6 == 5'd4) ? M_sheep : 0;
   assign M_sprite6 = (id6 == 5'd5) ? M_cow : 0;
   assign M_sprite6 = (id6 == 5'd6) ? M_hen : 0;
   assign M_sprite6 = (id6 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite6 = (id6 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite6 = (id6 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite6 = (id6 == 5'd10) ? M_score : 0;
   assign M_sprite6 = (id6 == 5'd11) ? M_one : 0;
   assign M_sprite6 = (id6 == 5'd12) ? M_two : 0;
   assign M_sprite6 = (id6 == 5'd13) ? M_three : 0;
   assign M_sprite6 = (id6 == 5'd14) ? M_four : 0;
   assign M_sprite6 = (id6 == 5'd15) ? M_five : 0;
   assign M_sprite6 = (id6 == 5'd16) ? M_six : 0;
   assign M_sprite6 = (id6 == 5'd17) ? M_seven : 0;
   assign M_sprite6 = (id6 == 5'd18) ? M_eight : 0;
   assign M_sprite6 = (id6 == 5'd19) ? M_nine : 0;
   assign M_sprite6 = (id6 == 5'd20) ? M_zero : 0;
   assign M_sprite6 = (id6 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite7 = (id7 == 5'd1) ? M_ship : 0;
   assign M_sprite7 = (id7 == 5'd2) ? M_pig : 0;
   assign M_sprite7 = (id7 == 5'd3) ? M_bee : 0;
   assign M_sprite7 = (id7 == 5'd4) ? M_sheep : 0;
   assign M_sprite7 = (id7 == 5'd5) ? M_cow : 0;
   assign M_sprite7 = (id7 == 5'd6) ? M_hen : 0;
   assign M_sprite7 = (id7 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite7 = (id7 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite7 = (id7 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite7 = (id7 == 5'd10) ? M_score : 0;
   assign M_sprite7 = (id7 == 5'd11) ? M_one : 0;
   assign M_sprite7 = (id7 == 5'd12) ? M_two : 0;
   assign M_sprite7 = (id7 == 5'd13) ? M_three : 0;
   assign M_sprite7 = (id7 == 5'd14) ? M_four : 0;
   assign M_sprite7 = (id7 == 5'd15) ? M_five : 0;
   assign M_sprite7 = (id7 == 5'd16) ? M_six : 0;
   assign M_sprite7 = (id7 == 5'd17) ? M_seven : 0;
   assign M_sprite7 = (id7 == 5'd18) ? M_eight : 0;
   assign M_sprite7 = (id7 == 5'd19) ? M_nine : 0;
   assign M_sprite7 = (id7 == 5'd20) ? M_zero : 0;
   assign M_sprite7 = (id7 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite8 = (id8 == 5'd1) ? M_ship : 0;
   assign M_sprite8 = (id8 == 5'd2) ? M_pig : 0;
   assign M_sprite8 = (id8 == 5'd3) ? M_bee : 0;
   assign M_sprite8 = (id8 == 5'd4) ? M_sheep : 0;
   assign M_sprite8 = (id8 == 5'd5) ? M_cow : 0;
   assign M_sprite8 = (id8 == 5'd6) ? M_hen : 0;
   assign M_sprite8 = (id8 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite8 = (id8 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite8 = (id8 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite8 = (id8 == 5'd10) ? M_score : 0;
   assign M_sprite8 = (id8 == 5'd11) ? M_one : 0;
   assign M_sprite8 = (id8 == 5'd12) ? M_two : 0;
   assign M_sprite8 = (id8 == 5'd13) ? M_three : 0;
   assign M_sprite8 = (id8 == 5'd14) ? M_four : 0;
   assign M_sprite8 = (id8 == 5'd15) ? M_five : 0;
   assign M_sprite8 = (id8 == 5'd16) ? M_six : 0;
   assign M_sprite8 = (id8 == 5'd17) ? M_seven : 0;
   assign M_sprite8 = (id8 == 5'd18) ? M_eight : 0;
   assign M_sprite8 = (id8 == 5'd19) ? M_nine : 0;
   assign M_sprite8 = (id8 == 5'd20) ? M_zero : 0;
   assign M_sprite8 = (id8 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite9 = (id9 == 5'd1) ? M_ship : 0;
   assign M_sprite9 = (id9 == 5'd2) ? M_pig : 0;
   assign M_sprite9 = (id9 == 5'd3) ? M_bee : 0;
   assign M_sprite9 = (id9 == 5'd4) ? M_sheep : 0;
   assign M_sprite9 = (id9 == 5'd5) ? M_cow : 0;
   assign M_sprite9 = (id9 == 5'd6) ? M_hen : 0;
   assign M_sprite9 = (id9 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite9 = (id9 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite9 = (id9 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite9 = (id9 == 5'd10) ? M_score : 0;
   assign M_sprite9 = (id9 == 5'd11) ? M_one : 0;
   assign M_sprite9 = (id9 == 5'd12) ? M_two : 0;
   assign M_sprite9 = (id9 == 5'd13) ? M_three : 0;
   assign M_sprite9 = (id9 == 5'd14) ? M_four : 0;
   assign M_sprite9 = (id9 == 5'd15) ? M_five : 0;
   assign M_sprite9 = (id9 == 5'd16) ? M_six : 0;
   assign M_sprite9 = (id9 == 5'd17) ? M_seven : 0;
   assign M_sprite9 = (id9 == 5'd18) ? M_eight : 0;
   assign M_sprite9 = (id9 == 5'd19) ? M_nine : 0;
   assign M_sprite9 = (id9 == 5'd20) ? M_zero : 0;
   assign M_sprite9 = (id9 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite10 = (id10 == 5'd1) ? M_ship : 0;
   assign M_sprite10 = (id10 == 5'd2) ? M_pig : 0;
   assign M_sprite10 = (id10 == 5'd3) ? M_bee : 0;
   assign M_sprite10 = (id10 == 5'd4) ? M_sheep : 0;
   assign M_sprite10 = (id10 == 5'd5) ? M_cow : 0;
   assign M_sprite10 = (id10 == 5'd6) ? M_hen : 0;
   assign M_sprite10 = (id10 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite10 = (id10 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite10 = (id10 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite10 = (id10 == 5'd10) ? M_score : 0;
   assign M_sprite10 = (id10 == 5'd11) ? M_one : 0;
   assign M_sprite10 = (id10 == 5'd12) ? M_two : 0;
   assign M_sprite10 = (id10 == 5'd13) ? M_three : 0;
   assign M_sprite10 = (id10 == 5'd14) ? M_four : 0;
   assign M_sprite10 = (id10 == 5'd15) ? M_five : 0;
   assign M_sprite10 = (id10 == 5'd16) ? M_six : 0;
   assign M_sprite10 = (id10 == 5'd17) ? M_seven : 0;
   assign M_sprite10 = (id10 == 5'd18) ? M_eight : 0;
   assign M_sprite10 = (id10 == 5'd19) ? M_nine : 0;
   assign M_sprite10 = (id10 == 5'd20) ? M_zero : 0;
   assign M_sprite10 = (id10 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite11 = (id11 == 5'd1) ? M_ship : 0;
   assign M_sprite11 = (id11 == 5'd2) ? M_pig : 0;
   assign M_sprite11 = (id11 == 5'd3) ? M_bee : 0;
   assign M_sprite11 = (id11 == 5'd4) ? M_sheep : 0;
   assign M_sprite11 = (id11 == 5'd5) ? M_cow : 0;
   assign M_sprite11 = (id11 == 5'd6) ? M_hen : 0;
   assign M_sprite11 = (id11 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite11 = (id11 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite11 = (id11 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite11 = (id11 == 5'd10) ? M_score : 0;
   assign M_sprite11 = (id11 == 5'd11) ? M_one : 0;
   assign M_sprite11 = (id11 == 5'd12) ? M_two : 0;
   assign M_sprite11 = (id11 == 5'd13) ? M_three : 0;
   assign M_sprite11 = (id11 == 5'd14) ? M_four : 0;
   assign M_sprite11 = (id11 == 5'd15) ? M_five : 0;
   assign M_sprite11 = (id11 == 5'd16) ? M_six : 0;
   assign M_sprite11 = (id11 == 5'd17) ? M_seven : 0;
   assign M_sprite11 = (id11 == 5'd18) ? M_eight : 0;
   assign M_sprite11 = (id11 == 5'd19) ? M_nine : 0;
   assign M_sprite11 = (id11 == 5'd20) ? M_zero : 0;
   assign M_sprite11 = (id11 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite12 = (id12 == 5'd1) ? M_ship : 0;
   assign M_sprite12 = (id12 == 5'd2) ? M_pig : 0;
   assign M_sprite12 = (id12 == 5'd3) ? M_bee : 0;
   assign M_sprite12 = (id12 == 5'd4) ? M_sheep : 0;
   assign M_sprite12 = (id12 == 5'd5) ? M_cow : 0;
   assign M_sprite12 = (id12 == 5'd6) ? M_hen : 0;
   assign M_sprite12 = (id12 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite12 = (id12 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite12 = (id12 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite12 = (id12 == 5'd10) ? M_score : 0;
   assign M_sprite12 = (id12 == 5'd11) ? M_one : 0;
   assign M_sprite12 = (id12 == 5'd12) ? M_two : 0;
   assign M_sprite12 = (id12 == 5'd13) ? M_three : 0;
   assign M_sprite12 = (id12 == 5'd14) ? M_four : 0;
   assign M_sprite12 = (id12 == 5'd15) ? M_five : 0;
   assign M_sprite12 = (id12 == 5'd16) ? M_six : 0;
   assign M_sprite12 = (id12 == 5'd17) ? M_seven : 0;
   assign M_sprite12 = (id12 == 5'd18) ? M_eight : 0;
   assign M_sprite12 = (id12 == 5'd19) ? M_nine : 0;
   assign M_sprite12 = (id12 == 5'd20) ? M_zero : 0;
   assign M_sprite12 = (id12 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite13 = (id13 == 5'd1) ? M_ship : 0;
   assign M_sprite13 = (id13 == 5'd2) ? M_pig : 0;
   assign M_sprite13 = (id13 == 5'd3) ? M_bee : 0;
   assign M_sprite13 = (id13 == 5'd4) ? M_sheep : 0;
   assign M_sprite13 = (id13 == 5'd5) ? M_cow : 0;
   assign M_sprite13 = (id13 == 5'd6) ? M_hen : 0;
   assign M_sprite13 = (id13 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite13 = (id13 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite13 = (id13 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite13 = (id13 == 5'd10) ? M_score : 0;
   assign M_sprite13 = (id13 == 5'd11) ? M_one : 0;
   assign M_sprite13 = (id13 == 5'd12) ? M_two : 0;
   assign M_sprite13 = (id13 == 5'd13) ? M_three : 0;
   assign M_sprite13 = (id13 == 5'd14) ? M_four : 0;
   assign M_sprite13 = (id13 == 5'd15) ? M_five : 0;
   assign M_sprite13 = (id13 == 5'd16) ? M_six : 0;
   assign M_sprite13 = (id13 == 5'd17) ? M_seven : 0;
   assign M_sprite13 = (id13 == 5'd18) ? M_eight : 0;
   assign M_sprite13 = (id13 == 5'd19) ? M_nine : 0;
   assign M_sprite13 = (id13 == 5'd20) ? M_zero : 0;
   assign M_sprite13 = (id13 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite14 = (id14 == 5'd1) ? M_ship : 0;
   assign M_sprite14 = (id14 == 5'd2) ? M_pig : 0;
   assign M_sprite14 = (id14 == 5'd3) ? M_bee : 0;
   assign M_sprite14 = (id14 == 5'd4) ? M_sheep : 0;
   assign M_sprite14 = (id14 == 5'd5) ? M_cow : 0;
   assign M_sprite14 = (id14 == 5'd6) ? M_hen : 0;
   assign M_sprite14 = (id14 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite14 = (id14 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite14 = (id14 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite14 = (id14 == 5'd10) ? M_score : 0;
   assign M_sprite14 = (id14 == 5'd11) ? M_one : 0;
   assign M_sprite14 = (id14 == 5'd12) ? M_two : 0;
   assign M_sprite14 = (id14 == 5'd13) ? M_three : 0;
   assign M_sprite14 = (id14 == 5'd14) ? M_four : 0;
   assign M_sprite14 = (id14 == 5'd15) ? M_five : 0;
   assign M_sprite14 = (id14 == 5'd16) ? M_six : 0;
   assign M_sprite14 = (id14 == 5'd17) ? M_seven : 0;
   assign M_sprite14 = (id14 == 5'd18) ? M_eight : 0;
   assign M_sprite14 = (id14 == 5'd19) ? M_nine : 0;
   assign M_sprite14 = (id14 == 5'd20) ? M_zero : 0;
   assign M_sprite14 = (id14 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite15 = (id15 == 5'd1) ? M_ship : 0;
   assign M_sprite15 = (id15 == 5'd2) ? M_pig : 0;
   assign M_sprite15 = (id15 == 5'd3) ? M_bee : 0;
   assign M_sprite15 = (id15 == 5'd4) ? M_sheep : 0;
   assign M_sprite15 = (id15 == 5'd5) ? M_cow : 0;
   assign M_sprite15 = (id15 == 5'd6) ? M_hen : 0;
   assign M_sprite15 = (id15 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite15 = (id15 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite15 = (id15 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite15 = (id15 == 5'd10) ? M_score : 0;
   assign M_sprite15 = (id15 == 5'd11) ? M_one : 0;
   assign M_sprite15 = (id15 == 5'd12) ? M_two : 0;
   assign M_sprite15 = (id15 == 5'd13) ? M_three : 0;
   assign M_sprite15 = (id15 == 5'd14) ? M_four : 0;
   assign M_sprite15 = (id15 == 5'd15) ? M_five : 0;
   assign M_sprite15 = (id15 == 5'd16) ? M_six : 0;
   assign M_sprite15 = (id15 == 5'd17) ? M_seven : 0;
   assign M_sprite15 = (id15 == 5'd18) ? M_eight : 0;
   assign M_sprite15 = (id15 == 5'd19) ? M_nine : 0;
   assign M_sprite15 = (id15 == 5'd20) ? M_zero : 0;
   assign M_sprite15 = (id15 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite16 = (id16 == 5'd1) ? M_ship : 0;
   assign M_sprite16 = (id16 == 5'd2) ? M_pig : 0;
   assign M_sprite16 = (id16 == 5'd3) ? M_bee : 0;
   assign M_sprite16 = (id16 == 5'd4) ? M_sheep : 0;
   assign M_sprite16 = (id16 == 5'd5) ? M_cow : 0;
   assign M_sprite16 = (id16 == 5'd6) ? M_hen : 0;
   assign M_sprite16 = (id16 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite16 = (id16 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite16 = (id16 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite16 = (id16 == 5'd10) ? M_score : 0;
   assign M_sprite16 = (id16 == 5'd11) ? M_one : 0;
   assign M_sprite16 = (id16 == 5'd12) ? M_two : 0;
   assign M_sprite16 = (id16 == 5'd13) ? M_three : 0;
   assign M_sprite16 = (id16 == 5'd14) ? M_four : 0;
   assign M_sprite16 = (id16 == 5'd15) ? M_five : 0;
   assign M_sprite16 = (id16 == 5'd16) ? M_six : 0;
   assign M_sprite16 = (id16 == 5'd17) ? M_seven : 0;
   assign M_sprite16 = (id16 == 5'd18) ? M_eight : 0;
   assign M_sprite16 = (id16 == 5'd19) ? M_nine : 0;
   assign M_sprite16 = (id16 == 5'd20) ? M_zero : 0;
   assign M_sprite16 = (id16 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite17 = (id17 == 5'd1) ? M_ship : 0;
   assign M_sprite17 = (id17 == 5'd2) ? M_pig : 0;
   assign M_sprite17 = (id17 == 5'd3) ? M_bee : 0;
   assign M_sprite17 = (id17 == 5'd4) ? M_sheep : 0;
   assign M_sprite17 = (id17 == 5'd5) ? M_cow : 0;
   assign M_sprite17 = (id17 == 5'd6) ? M_hen : 0;
   assign M_sprite17 = (id17 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite17 = (id17 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite17 = (id17 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite17 = (id17 == 5'd10) ? M_score : 0;
   assign M_sprite17 = (id17 == 5'd11) ? M_one : 0;
   assign M_sprite17 = (id17 == 5'd12) ? M_two : 0;
   assign M_sprite17 = (id17 == 5'd13) ? M_three : 0;
   assign M_sprite17 = (id17 == 5'd14) ? M_four : 0;
   assign M_sprite17 = (id17 == 5'd15) ? M_five : 0;
   assign M_sprite17 = (id17 == 5'd16) ? M_six : 0;
   assign M_sprite17 = (id17 == 5'd17) ? M_seven : 0;
   assign M_sprite17 = (id17 == 5'd18) ? M_eight : 0;
   assign M_sprite17 = (id17 == 5'd19) ? M_nine : 0;
   assign M_sprite17 = (id17 == 5'd20) ? M_zero : 0;
   assign M_sprite17 = (id17 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite18 = (id18 == 5'd1) ? M_ship : 0;
   assign M_sprite18 = (id18 == 5'd2) ? M_pig : 0;
   assign M_sprite18 = (id18 == 5'd3) ? M_bee : 0;
   assign M_sprite18 = (id18 == 5'd4) ? M_sheep : 0;
   assign M_sprite18 = (id18 == 5'd5) ? M_cow : 0;
   assign M_sprite18 = (id18 == 5'd6) ? M_hen : 0;
   assign M_sprite18 = (id18 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite18 = (id18 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite18 = (id18 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite18 = (id18 == 5'd10) ? M_score : 0;
   assign M_sprite18 = (id18 == 5'd11) ? M_one : 0;
   assign M_sprite18 = (id18 == 5'd12) ? M_two : 0;
   assign M_sprite18 = (id18 == 5'd13) ? M_three : 0;
   assign M_sprite18 = (id18 == 5'd14) ? M_four : 0;
   assign M_sprite18 = (id18 == 5'd15) ? M_five : 0;
   assign M_sprite18 = (id18 == 5'd16) ? M_six : 0;
   assign M_sprite18 = (id18 == 5'd17) ? M_seven : 0;
   assign M_sprite18 = (id18 == 5'd18) ? M_eight : 0;
   assign M_sprite18 = (id18 == 5'd19) ? M_nine : 0;
   assign M_sprite18 = (id18 == 5'd20) ? M_zero : 0;
   assign M_sprite18 = (id18 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite19 = (id19 == 5'd1) ? M_ship : 0;
   assign M_sprite19 = (id19 == 5'd2) ? M_pig : 0;
   assign M_sprite19 = (id19 == 5'd3) ? M_bee : 0;
   assign M_sprite19 = (id19 == 5'd4) ? M_sheep : 0;
   assign M_sprite19 = (id19 == 5'd5) ? M_cow : 0;
   assign M_sprite19 = (id19 == 5'd6) ? M_hen : 0;
   assign M_sprite19 = (id19 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite19 = (id19 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite19 = (id19 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite19 = (id19 == 5'd10) ? M_score : 0;
   assign M_sprite19 = (id19 == 5'd11) ? M_one : 0;
   assign M_sprite19 = (id19 == 5'd12) ? M_two : 0;
   assign M_sprite19 = (id19 == 5'd13) ? M_three : 0;
   assign M_sprite19 = (id19 == 5'd14) ? M_four : 0;
   assign M_sprite19 = (id19 == 5'd15) ? M_five : 0;
   assign M_sprite19 = (id19 == 5'd16) ? M_six : 0;
   assign M_sprite19 = (id19 == 5'd17) ? M_seven : 0;
   assign M_sprite19 = (id19 == 5'd18) ? M_eight : 0;
   assign M_sprite19 = (id19 == 5'd19) ? M_nine : 0;
   assign M_sprite19 = (id19 == 5'd20) ? M_zero : 0;
   assign M_sprite19 = (id19 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite20 = (id20 == 5'd1) ? M_ship : 0;
   assign M_sprite20 = (id20 == 5'd2) ? M_pig : 0;
   assign M_sprite20 = (id20 == 5'd3) ? M_bee : 0;
   assign M_sprite20 = (id20 == 5'd4) ? M_sheep : 0;
   assign M_sprite20 = (id20 == 5'd5) ? M_cow : 0;
   assign M_sprite20 = (id20 == 5'd6) ? M_hen : 0;
   assign M_sprite20 = (id20 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite20 = (id20 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite20 = (id20 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite20 = (id20 == 5'd10) ? M_score : 0;
   assign M_sprite20 = (id20 == 5'd11) ? M_one : 0;
   assign M_sprite20 = (id20 == 5'd12) ? M_two : 0;
   assign M_sprite20 = (id20 == 5'd13) ? M_three : 0;
   assign M_sprite20 = (id20 == 5'd14) ? M_four : 0;
   assign M_sprite20 = (id20 == 5'd15) ? M_five : 0;
   assign M_sprite20 = (id20 == 5'd16) ? M_six : 0;
   assign M_sprite20 = (id20 == 5'd17) ? M_seven : 0;
   assign M_sprite20 = (id20 == 5'd18) ? M_eight : 0;
   assign M_sprite20 = (id20 == 5'd19) ? M_nine : 0;
   assign M_sprite20 = (id20 == 5'd20) ? M_zero : 0;
   assign M_sprite20 = (id20 == 5'd21) ? M_bullet : 0;
   
   assign M_sprite21 = (id21 == 5'd1) ? M_ship : 0;
   assign M_sprite21 = (id21 == 5'd2) ? M_pig : 0;
   assign M_sprite21 = (id21 == 5'd3) ? M_bee : 0;
   assign M_sprite21 = (id21 == 5'd4) ? M_sheep : 0;
   assign M_sprite21 = (id21 == 5'd5) ? M_cow : 0;
   assign M_sprite21 = (id21 == 5'd6) ? M_hen : 0;
   assign M_sprite21 = (id21 == 5'd7) ? M_mcdonald : 0;
   assign M_sprite21 = (id21 == 5'd8) ? M_h_eskimo : 0;
   assign M_sprite21 = (id21 == 5'd9) ? M_s_eskimo : 0;
   assign M_sprite21 = (id21 == 5'd10) ? M_score : 0;
   assign M_sprite21 = (id21 == 5'd11) ? M_one : 0;
   assign M_sprite21 = (id21 == 5'd12) ? M_two : 0;
   assign M_sprite21 = (id21 == 5'd13) ? M_three : 0;
   assign M_sprite21 = (id21 == 5'd14) ? M_four : 0;
   assign M_sprite21 = (id21 == 5'd15) ? M_five : 0;
   assign M_sprite21 = (id21 == 5'd16) ? M_six : 0;
   assign M_sprite21 = (id21 == 5'd17) ? M_seven : 0;
   assign M_sprite21 = (id21 == 5'd18) ? M_eight : 0;
   assign M_sprite21 = (id21 == 5'd19) ? M_nine : 0;
   assign M_sprite21 = (id20 == 5'd20) ? M_zero : 0;
   assign M_sprite21 = (id21 == 5'd21) ? M_bullet : 0;
   

   ship mn(.clock(VGA_CLK), .address(addr_ship), .q(M_ship));
   pig mn(.clock(VGA_CLK), .address(addr_pig), .q(M_pig));
   bee mn(.clock(VGA_CLK), .address(addr_bee), .q(M_bee));
   sheep mn(.clock(VGA_CLK), .address(addr_sheep), .q(M_sheep));
   cow mn(.clock(VGA_CLK), .address(addr_cow), .q(M_cow));
   hen mn(.clock(VGA_CLK), .address(addr_hen), .q(M_hen));
   mcdonald mn(.clock(VGA_CLK), .address(addr_mcdonald), .q(M_mcdonald));
   h_eskimo mn(.clock(VGA_CLK), .address(addr_h_eskimo), .q(M_h_eskimo));
   s_eskimo mn(.clock(VGA_CLK), .address(addr_s_eskimo), .q(M_s_eskimo));
   score mn(.clock(VGA_CLK), .address(addr_score), .q(M_score));
   one mn(.clock(VGA_CLK), .address(addr_one), .q(M_one));
   two mn(.clock(VGA_CLK), .address(addr_two), .q(M_two));
   three mn(.clock(VGA_CLK), .address(addr_three), .q(M_three));
   four mn(.clock(VGA_CLK), .address(addr_four), .q(M_four));
   five mn(.clock(VGA_CLK), .address(addr_five), .q(M_five));
   six mn(.clock(VGA_CLK), .address(addr_six), .q(M_six));
   seven mn(.clock(VGA_CLK), .address(addr_seven), .q(M_seven));
   eight mn(.clock(VGA_CLK), .address(addr_eight), .q(M_eight));
   nine mn(.clock(VGA_CLK), .address(addr_nine), .q(M_nine));
   zero mn(.clock(VGA_CLK), .address(addr_zero), .q(M_zero));
   bullet mn(.clock(VGA_CLK), .address(addr_bullet), .q(M_bullet));

   

   VGA_LED_Emulator led_emulator(.clk50(clk), .*);
   Sprite_Controller sprite_controller(.clk(VGA_CLK), .sprite1(gl_array[0]), .*);

endmodule
